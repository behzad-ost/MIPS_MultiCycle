library verilog;
use verilog.vl_types.all;
entity CPU_test is
end CPU_test;
